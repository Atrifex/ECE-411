library verilog;
use verilog.vl_types.all;
entity way_sv_unit is
end way_sv_unit;
