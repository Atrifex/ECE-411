library verilog;
use verilog.vl_types.all;
entity cache_writelogic_sv_unit is
end cache_writelogic_sv_unit;
